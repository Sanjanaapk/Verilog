module not2(
 input x,
 output f);
 assign f = ~x;
 endmodule